module rotright_gate(
	input wire [31:0] A,
	input wire [4:0] B, 
	output wire [31:0] out
);

reg [31:0] C;

always@(*) begin
	case(B)
		5'd31: C <= {A[30:0], A[31]};
		5'd30: C <= {A[29:0], A[31:30]};
		5'd29: C <= {A[28:0], A[31:29]};
		5'd28: C <= {A[27:0], A[31:28]};
		5'd27: C <= {A[26:0], A[31:27]};
		5'd26: C <= {A[25:0], A[31:26]};
		5'd25: C <= {A[24:0], A[31:25]};
		5'd24: C <= {A[23:0], A[31:24]};
		5'd23: C <= {A[22:0], A[31:23]};
		5'd22: C <= {A[21:0], A[31:22]};
		5'd21: C <= {A[20:0], A[31:21]};
		5'd20: C <= {A[19:0], A[31:20]};
		5'd19: C <= {A[18:0], A[31:19]};
		5'd18: C <= {A[17:0], A[31:18]};
		5'd17: C <= {A[16:0], A[31:17]};
		5'd16: C <= {A[15:0], A[31:16]};
		5'd15: C <= {A[14:0], A[31:15]};
		5'd14: C <= {A[13:0], A[31:14]};
		5'd13: C <= {A[12:0], A[31:13]};
		5'd12: C <= {A[11:0], A[31:12]};
		5'd11: C <= {A[10:0], A[31:11]};
		5'd10: C <= {A[9:0], A[31:10]};
		5'd9: C <= {A[8:0], A[31:9]};
		5'd8: C <= {A[7:0], A[31:8]};
		5'd7: C <= {A[6:0], A[31:7]};
		5'd6: C <= {A[5:0], A[31:6]};
		5'd5: C <= {A[4:0], A[31:5]};
		5'd4: C <= {A[3:0], A[31:4]};
		5'd3: C <= {A[2:0], A[31:3]};
		5'd2:	C <= {A[1:0], A[31:2]};
		5'd1:	C <= {A[0], A[31:1]};
		default: C <= A;
	endcase
end  
assign out = C;
endmodule 