module or_gate(
	input wire [31:0] A, B, 
	output wire [31:0] C
);

assign C = A | B;
endmodule 